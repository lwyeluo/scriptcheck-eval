https://www.google.com.sv/
